----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
--
library altera;
use altera.altera_primitives_components.all;
library work;
use work.global_def_package.all;
use work.xge_package.all;
use work.test_package.all;
use work.s5_source_probe_package.all;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
entity top is
	generic
	(
		DEF_TB_ROLE											: t_tb_role := SLAVE
	);
	port
	(
		-- CLOCK
		i_clk_50_B3B										: in std_logic := '0';
		i_clk_50_B3D										: in std_logic := '0';
		i_clk_50_B4A										: in std_logic := '0';
		i_clk_50_B4D										: in std_logic := '0';
		i_clk_50_B7A										: in std_logic := '0';
		i_clk_50_B7D										: in std_logic := '0';
		i_clk_50_B8A										: in std_logic := '0';
		i_clk_50_B8D										: in std_logic := '0';
		-- LED x 10
		o_LED												: out std_logic_vector(3 downto 0) := (others => '0');
		o_LED_BRACKET										: out std_logic_vector(3 downto 0) := (others => '0');
		o_LED_RJ45_L										: out std_logic := '0';
		o_LED_RJ45_R										: out std_logic := '0';
		-- BUTTON x 4 and CPU_RESET_n
		i_BUTTONS											: in std_logic_vector(3 downto 0) := (others => '0');
		i_CPU_RESET_n										: in std_logic := '0';
		-- SFP+ A
		i_SFPA_LOS											: in std_logic := '0';
		i_SFPA_MOD0_PRSNT_n									: in std_logic := '0';
		o_SFPA_MOD1_SCL										: out std_logic := '0';
		io_SFPA_MOD2_SDA									: inout std_logic := '0';
		o_SFPA_RATESEL										: out std_logic_vector(1 downto 0) := (others => '0');
		i_SFPA_RX_p											: in std_logic := '0';
		o_SFPA_TX_p											: out std_logic := '0';
		o_SFPA_TXDISABLE									: out std_logic := '0';
		i_SFPA_TXFAULT										: in std_logic := '0';
		-- SFP+ B
		i_SFPB_LOS											: in std_logic := '0';
		i_SFPB_MOD0_PRSNT_n									: in std_logic := '0';
		o_SFPB_MOD1_SCL										: out std_logic := '0';
		io_SFPB_MOD2_SDA									: inout std_logic := '0';
		o_SFPB_RATESEL										: out std_logic_vector(1 downto 0) := (others => '0');
		i_SFPB_RX_p											: in std_logic := '0';
		o_SFPB_TX_p											: out std_logic := '0';
		o_SFPB_TXDISABLE									: out std_logic := '0';
		i_SFPB_TXFAULT										: in std_logic := '0';
		-- SFP+ C
		i_SFPC_LOS											: in std_logic := '0';
		i_SFPC_MOD0_PRSNT_n									: in std_logic := '0';
		o_SFPC_MOD1_SCL										: out std_logic := '0';
		io_SFPC_MOD2_SDA									: inout std_logic := '0';
		o_SFPC_RATESEL										: out std_logic_vector(1 downto 0) := (others => '0');
		i_SFPC_RX_p											: in std_logic := '0';
		o_SFPC_TX_p											: out std_logic := '0';
		o_SFPC_TXDISABLE									: out std_logic := '0';
		i_SFPC_TXFAULT										: in std_logic := '0';
		-- SFP+ D
		i_SFPD_LOS											: in std_logic := '0';
		i_SFPD_MOD0_PRSNT_n									: in std_logic := '0';
		o_SFPD_MOD1_SCL										: out std_logic := '0';
		io_SFPD_MOD2_SDA									: inout std_logic := '0';
		o_SFPD_RATESEL										: out std_logic_vector(1 downto 0) := (others => '0');
		i_SFPD_RX_p											: in std_logic := '0';
		o_SFPD_TX_p											: out std_logic := '0';
		o_SFPD_TXDISABLE									: out std_logic := '0';
		i_SFPD_TXFAULT										: in std_logic := '0';
		-- SFP+ 10G Referece Clock (generated by the Programmalbe Oscillator Si570)
		i_SFP_REFCLK_p										: in std_logic := '0';
		-- Programmalbe Oscillator SI570
		o_CLOCK_SCL											: out std_logic := '0';
		io_CLOCK_SDA										: inout std_logic := '0';
		-- Fan
		io_FAN_CTRL											: inout std_logic := '0';
		-- Temperature
		o_TEMP_CLK											: out std_logic := '0';
		io_TEMP_DATA										: inout std_logic := '0';
		i_TEMP_INT_n										: in std_logic := '0';
		i_TEMP_OVERT_n										: in std_logic := '0'
	);
end entity;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
architecture rtl of top is
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
component xge_main is
	generic
	(
		DEF_TB_ROLE											: t_tb_role := SLAVE
	);
	port
	(
		i_clk_50											: in std_logic := '0';
		i_reset												: in std_logic := '0';
		--
		i_xge_tx_pll_refclk									: in std_logic := '0';
		i_xge_rx_cdr_refclk									: in std_logic := '0';
		--
		o_xge_N_tx_serial_data								: out std_logic_vector(C_SFP_N_CHANNEL-1 downto 0) := (others => '0');
		i_xge_N_rx_serial_data								: in std_logic_vector(C_SFP_N_CHANNEL-1 downto 0) := (others => '0');
		--
		i_rcd_source_probe									: in t_rcd_s5_source_probe := ci_t_rcd_s5_source_probe;
		i_rcd_temperature									: in t_rcd_temperature := ci_t_rcd_temperature
	);
end component;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
component si570_controller
	port
	(
		iCLK												: in std_logic := '0';										-- system clock 50mhz 
		iRST_n												: in std_logic := '0';										-- system reset;
		iStart												: in std_logic := '0';
		iFREQ_MODE											: in std_logic_vector(2 downto 0) := (others => '0');
		I2C_CLK												: out std_logic := '0';
		I2C_DATA											: inout std_logic := '0';
		oController_Ready									: out std_logic := '0'
	);
end component;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
component cmp_s5_pll_644 is
	port
	(
		refclk												: in std_logic := '0';
		rst													: in std_logic := '0';
		outclk_0 											: out std_logic;
		locked												: out std_logic
	);
end component;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
component s5_source_probe is
	port
	(
		i_clk												: in std_logic := '0';
		o_rcd												: out t_rcd_s5_source_probe := ci_t_rcd_s5_source_probe
	);
end component;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
component s5_temperature is
	port
	(
		i_clk								: in std_logic := '0';										-- 50МГц
		o_TEMP_CLK							: out std_logic := '1';										-- i2c
		io_TEMP_DATA						: inout std_logic := '1';									-- i2c
		o_TempByte							: out std_logic_vector(7 downto 0) := (others => '0');		-- результирующее прочитанное слово
		--
		o_TempByte_L_valid					: out std_logic := '0';										-- 
		o_TempByte_L						: out std_logic_vector(7 downto 0) := (others => '0');		-- 
		o_TempByte_R_valid					: out std_logic := '0';										-- 
		o_TempByte_R						: out std_logic_vector(7 downto 0) := (others => '0');		-- 
		o_TempByte_MAN_ID_valid				: out std_logic := '0';										-- 
		o_TempByte_MAN_ID					: out std_logic_vector(7 downto 0) := (others => '0');		-- 
		o_TempByte_DEV_ID_valid				: out std_logic := '0';										-- 
		o_TempByte_DEV_ID					: out std_logic_vector(7 downto 0) := (others => '0')		-- 
	);
end component;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
constant CT_ANTI_SHATTER									: integer := 50000;
--
signal cpu_reset_2w_clk50									: std_logic := '0';
signal cpu_reset_2w_clk50_last								: std_logic := '0';
--
signal cpu_reset_n_z0										: std_logic := '0';
signal cpu_reset_n_z1										: std_logic := '0';
signal cpu_reset_n_z1_last									: std_logic := '0';
signal cpu_reset_n_cnt										: integer range 0 to CT_ANTI_SHATTER + 10 := 0;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
constant CT_SI570_FREQ_MODE									: std_logic_vector(2 downto 0) := "110";
constant CT_SI570_TIME_CMD_RESET							: integer := 100;
constant CT_SI570_TIME_CMD_START							: integer := 200;
constant CT_SI570_CMD_INTERVAL								: integer := 50;
signal si570_reset											: std_logic := '0';
signal si570_reset_n										: std_logic := '0';
signal si570_start											: std_logic := '0';
signal si570_cnt											: integer range 0 to CT_SI570_TIME_CMD_START + CT_SI570_CMD_INTERVAL + 10 := 0;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
signal xge_reset											: std_logic := '0';
signal xge_N_tx_serial_data									: std_logic_vector(C_SFP_N_CHANNEL-1 downto 0) := (others => '0');
signal xge_N_rx_serial_data									: std_logic_vector(C_SFP_N_CHANNEL-1 downto 0) := (others => '0');
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
signal s5_source_probe_o_rcd								: t_rcd_s5_source_probe := ci_t_rcd_s5_source_probe;
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
signal cmp_s5_pll_644_i_rst									: std_logic := '0';
signal cmp_s5_pll_644_o_clk_50								: std_logic := '0';
signal cmp_s5_pll_644_o_locked								: std_logic := '0';
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
signal fan_init_f											: std_logic := '0';
signal fan_turn_on_prev										: std_logic := '0';
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
signal rcd_s5_temperature									: t_rcd_temperature := ci_t_rcd_temperature;
signal s5_temperature_o_TempByte							: std_logic_vector(7 downto 0) := (others => '0');
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
signal LEDS													: std_logic_vector(3 downto 0) := (others => '0');
signal led0_cnt												: std_logic_vector(31 downto 0) := (others => '0');
signal led1_cnt												: std_logic_vector(31 downto 0) := (others => '0');
----------------------------------------------------------------------------------------------------------------------------------------------------------------------------
begin
	
	
	--======================================================================================================================================================================
	-- 10G ethernet (xge)
	--======================================================================================================================================================================
	xge_reset												<= cpu_reset_2w_clk50;
	---------------------------------------------
	gen_sfpa_0: if (C_SFP_N_CHANNEL > 0) generate
		o_SFPA_TX_p											<= xge_N_tx_serial_data(0);
		xge_N_rx_serial_data(0)								<= i_SFPA_RX_p;
	end generate;
	---------------------------------------------
	gen_sfpb_0: if (C_SFP_N_CHANNEL > 1) generate
		o_SFPB_TX_p											<= xge_N_tx_serial_data(1);
		xge_N_rx_serial_data(1)								<= i_SFPB_RX_p;
	end generate;
	gen_sfpb_1: if (C_SFP_N_CHANNEL < 2) generate
		o_SFPB_TX_p											<= i_SFPB_RX_p;
	end generate;
	---------------------------------------------
	gen_sfpc_0: if (C_SFP_N_CHANNEL > 2) generate
		o_SFPC_TX_p											<= xge_N_tx_serial_data(2);
		xge_N_rx_serial_data(2)								<= i_SFPC_RX_p;
	end generate;
	gen_sfpc_1: if (C_SFP_N_CHANNEL < 3) generate
		o_SFPC_TX_p											<= i_SFPC_RX_p;
	end generate;
	---------------------------------------------
	gen_sfpd_0: if (C_SFP_N_CHANNEL > 3) generate
		o_SFPD_TX_p											<= xge_N_tx_serial_data(3);
		xge_N_rx_serial_data(3)								<= i_SFPD_RX_p;
	end generate;
	gen_sfpd_1: if (C_SFP_N_CHANNEL < 4) generate
		o_SFPD_TX_p											<= i_SFPD_RX_p;
	end generate;
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	xge_main_x : xge_main
	generic map
	(
		DEF_TB_ROLE											=> DEF_TB_ROLE
	)
	port map
	(
		i_clk_50											=> i_clk_50_B3B,
		i_reset												=> xge_reset,
		--
		i_xge_tx_pll_refclk									=> i_SFP_REFCLK_p,		-- 644.53125 MHz
		i_xge_rx_cdr_refclk									=> i_SFP_REFCLK_p,		-- 644.53125 MHz
		--
		o_xge_N_tx_serial_data								=> xge_N_tx_serial_data,
		i_xge_N_rx_serial_data								=> xge_N_rx_serial_data,
		--
		i_rcd_source_probe									=> s5_source_probe_o_rcd,
		i_rcd_temperature									=> rcd_s5_temperature
	);
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	process(i_clk_50_B3B)
	begin
		if (rising_edge(i_clk_50_B3B)) then
			if (s5_source_probe_o_rcd.sfp.valid = '1') then
				o_SFPA_RATESEL								<= s5_source_probe_o_rcd.sfp.RATESEL;
				o_SFPA_TXDISABLE							<= s5_source_probe_o_rcd.sfp.TXDISABLE;
				o_SFPB_RATESEL								<= s5_source_probe_o_rcd.sfp.RATESEL;
				o_SFPB_TXDISABLE							<= s5_source_probe_o_rcd.sfp.TXDISABLE;
				o_SFPC_RATESEL								<= s5_source_probe_o_rcd.sfp.RATESEL;
				o_SFPC_TXDISABLE							<= s5_source_probe_o_rcd.sfp.TXDISABLE;
				o_SFPD_RATESEL								<= s5_source_probe_o_rcd.sfp.RATESEL;
				o_SFPD_TXDISABLE							<= s5_source_probe_o_rcd.sfp.TXDISABLE;
			else
				o_SFPA_RATESEL								<= (others => '0');
				o_SFPA_TXDISABLE							<= '0';
				o_SFPB_RATESEL								<= (others => '0');
				o_SFPB_TXDISABLE							<= '0';
				o_SFPC_RATESEL								<= (others => '0');
				o_SFPC_TXDISABLE							<= '0';
				o_SFPD_RATESEL								<= (others => '0');
				o_SFPD_TXDISABLE							<= '0';
			end if;
		end if;
	end process;
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	
	--======================================================================================================================================================================
	-- антидребезг i_CPU_RESET_n
	--======================================================================================================================================================================
	-- выходной сигнал:
	-- cpu_reset_2w_clk50
	process(i_clk_50_B3B)
	begin
		if (rising_edge(i_clk_50_B3B)) then
			cpu_reset_2w_clk50_last							<= cpu_reset_2w_clk50;
			if (cpu_reset_2w_clk50_last = '1') then
				cpu_reset_2w_clk50							<= '0';
			end if;
			--
			cpu_reset_n_z0									<= i_CPU_RESET_n;
			cpu_reset_n_z1									<= cpu_reset_n_z0;
			cpu_reset_n_z1_last								<= cpu_reset_n_z1;
			--
			if (cpu_reset_n_z1 = '0' AND cpu_reset_n_z1_last = '1' AND cpu_reset_n_cnt = 0) then
				cpu_reset_2w_clk50							<= '1';
				cpu_reset_n_cnt								<= 1;
			end if;
			if (cpu_reset_n_cnt > 0) then
				cpu_reset_n_cnt								<= cpu_reset_n_cnt + 1;
			end if;
			if (cpu_reset_n_cnt > CT_ANTI_SHATTER) then
				cpu_reset_n_cnt								<= 0;
			end if;
		end if;
	end process;
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	
	
	--======================================================================================================================================================================
	-- Configure SI570 as 644.5312 MHz
	--======================================================================================================================================================================
	process(i_clk_50_B3B)
	begin
		if (rising_edge(i_clk_50_B3B)) then
			if (cpu_reset_2w_clk50 = '1') then
				si570_reset									<= '0';
				si570_start									<= '0';
				si570_cnt									<= 0;
			else
				if (si570_cnt < CT_SI570_TIME_CMD_RESET) then
					si570_reset								<= '0';
					si570_start								<= '0';
					si570_cnt								<= si570_cnt + 1;
				elsif (si570_cnt >= CT_SI570_TIME_CMD_RESET AND si570_cnt < CT_SI570_TIME_CMD_RESET + CT_SI570_CMD_INTERVAL) then
					si570_reset								<= '1';
					si570_start								<= '0';
					si570_cnt								<= si570_cnt + 1;
				elsif (si570_cnt < CT_SI570_TIME_CMD_START) then
					si570_reset								<= '0';
					si570_start								<= '0';
					si570_cnt								<= si570_cnt + 1;
				elsif (si570_cnt >= CT_SI570_TIME_CMD_START AND si570_cnt < CT_SI570_TIME_CMD_START + CT_SI570_CMD_INTERVAL) then
					si570_reset								<= '0';
					si570_start								<= '1';
					si570_cnt								<= si570_cnt + 1;
				else
					si570_reset								<= '0';
					si570_start								<= '0';
				end if;
			end if;
		end if;
	end process;
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	si570_reset_n											<= not si570_reset;
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	si570_controller_x : si570_controller
	port map
	(
		iCLK												=> i_clk_50_B3B,		-- system clock 50mhz 
		iRST_n												=> si570_reset_n,		-- system reset;
		iStart												=> si570_start,
		iFREQ_MODE											=> CT_SI570_FREQ_MODE,
		I2C_CLK												=> o_CLOCK_SCL,
		I2C_DATA											=> io_CLOCK_SDA,
		oController_Ready									=> open
	);
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	
	
	--======================================================================================================================================================================
	-- Source Probe (Virtual Buttons)
	--======================================================================================================================================================================
	s5_source_probe_x : s5_source_probe
	port map
	(
		i_clk												=> i_clk_50_B3B,		-- system clock 50mhz 
		o_rcd												=> s5_source_probe_o_rcd
	);
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	
	
	--======================================================================================================================================================================
	-- Source Probe (Virtual Buttons)
	--======================================================================================================================================================================
	cmp_s5_pll_644_x : cmp_s5_pll_644
	port map
	(
		refclk												=> i_SFP_REFCLK_p,
		rst													=> cmp_s5_pll_644_i_rst,
		outclk_0 											=> cmp_s5_pll_644_o_clk_50,
		locked												=> cmp_s5_pll_644_o_locked
	);
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	
	
	--======================================================================================================================================================================
	-- LEDS
	--======================================================================================================================================================================
	o_LED(0)												<= LEDS(0);
	o_LED(1)												<= LEDS(1);
	o_LED(2)												<= LEDS(2);
	o_LED(3)												<= i_BUTTONS(3);
	--
	process(i_clk_50_B3B)
	begin
		if (rising_edge(i_clk_50_B3B)) then
			led0_cnt										<= led0_cnt + 1;
			LEDS(0)											<= led0_cnt(25);
		end if;	
	end process;
	--
	process(cmp_s5_pll_644_o_clk_50)
	begin
		if (rising_edge(cmp_s5_pll_644_o_clk_50)) then
			led1_cnt										<= led1_cnt + 1;
			LEDS(1)											<= led1_cnt(24);
		end if;	
	end process;
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	
	
	--======================================================================================================================================================================
	-- FAN
	--======================================================================================================================================================================
	process(i_clk_50_B3B)
	begin
		if (rising_edge(i_clk_50_B3B)) then
			if (fan_init_f = '0') then
				fan_init_f									<= '1';
				io_FAN_CTRL									<= '1';
			end if;
			--
			fan_turn_on_prev								<= s5_source_probe_o_rcd.main.fan_turn_on;
			if (s5_source_probe_o_rcd.main.fan_turn_on /= fan_turn_on_prev) then
				io_FAN_CTRL									<= s5_source_probe_o_rcd.main.fan_turn_on;
			end if;
		end if;	
	end process;
	------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	
	--======================================================================================================================================================================
	-- TTemperature MAX1619
	--======================================================================================================================================================================
	s5_temperature_x : s5_temperature
	port map
	(
		i_clk												=> i_clk_50_B3B,
		o_TEMP_CLK											=> o_TEMP_CLK,
		io_TEMP_DATA										=> io_TEMP_DATA,
		o_TempByte											=> s5_temperature_o_TempByte,
		--
		o_TempByte_L_valid									=> rcd_s5_temperature.T_L_valid,
		o_TempByte_L										=> rcd_s5_temperature.T_L,
		o_TempByte_R_valid									=> rcd_s5_temperature.T_R_valid,
		o_TempByte_R										=> rcd_s5_temperature.T_R,
		o_TempByte_MAN_ID_valid								=> rcd_s5_temperature.MAN_ID_valid,
		o_TempByte_MAN_ID									=> rcd_s5_temperature.MAN_ID,
		o_TempByte_DEV_ID_valid								=> rcd_s5_temperature.DEV_ID_valid,
		o_TempByte_DEV_ID									=> rcd_s5_temperature.DEV_ID
	);
	
end rtl;
